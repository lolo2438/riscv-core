library ieee;
use ieee.math_real.all;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_textio.all;
use std.textio.all;

entity XXX_tb is
end entity XXX_tb;

architecture test_bench of XXX_tb is

-- UUT SIGNALS



-- OTHER SIGNALS


begin




end architecture test_bench;
